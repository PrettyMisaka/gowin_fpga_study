module my_top(

);



endmodule