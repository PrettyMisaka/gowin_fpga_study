`ifndef __INOUT_H__
`define __INOUT_H__

interface inout_interface(
    input mdio_i,
    output logic mdio_o,
    output logic out_en
);
endinterface 

`endif
