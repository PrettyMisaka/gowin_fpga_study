`ifndef __CONFIG_H__
`define __CONFIG_H__

`include "rmii.svh"
`include "udp_interface.svh"
`include "cam_interface.svh"
`include "ddr3_interface.svh"

`endif