//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-5
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Sat Nov 04 19:29:56 2023

module Gowin_DPB_128_2048 (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [127:0] douta;
output [127:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [10:0] ada;
input [127:0] dina;
input [10:0] adb;
input [127:0] dinb;

wire [15:0] dpb_inst_0_douta;
wire [15:0] dpb_inst_0_doutb;
wire [15:0] dpb_inst_1_douta;
wire [15:0] dpb_inst_1_doutb;
wire [31:16] dpb_inst_2_douta;
wire [31:16] dpb_inst_2_doutb;
wire [31:16] dpb_inst_3_douta;
wire [31:16] dpb_inst_3_doutb;
wire [47:32] dpb_inst_4_douta;
wire [47:32] dpb_inst_4_doutb;
wire [47:32] dpb_inst_5_douta;
wire [47:32] dpb_inst_5_doutb;
wire [63:48] dpb_inst_6_douta;
wire [63:48] dpb_inst_6_doutb;
wire [63:48] dpb_inst_7_douta;
wire [63:48] dpb_inst_7_doutb;
wire [79:64] dpb_inst_8_douta;
wire [79:64] dpb_inst_8_doutb;
wire [79:64] dpb_inst_9_douta;
wire [79:64] dpb_inst_9_doutb;
wire [95:80] dpb_inst_10_douta;
wire [95:80] dpb_inst_10_doutb;
wire [95:80] dpb_inst_11_douta;
wire [95:80] dpb_inst_11_doutb;
wire [111:96] dpb_inst_12_douta;
wire [111:96] dpb_inst_12_doutb;
wire [111:96] dpb_inst_13_douta;
wire [111:96] dpb_inst_13_doutb;
wire [127:112] dpb_inst_14_douta;
wire [127:112] dpb_inst_14_doutb;
wire [127:112] dpb_inst_15_douta;
wire [127:112] dpb_inst_15_doutb;
wire dff_q_0;
wire dff_q_1;
wire cea_w;
wire ceb_w;
wire gw_vcc;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA(dpb_inst_0_douta[15:0]),
    .DOB(dpb_inst_0_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 16;
defparam dpb_inst_0.BIT_WIDTH_1 = 16;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";

DPB dpb_inst_1 (
    .DOA(dpb_inst_1_douta[15:0]),
    .DOB(dpb_inst_1_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_1.READ_MODE0 = 1'b0;
defparam dpb_inst_1.READ_MODE1 = 1'b0;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 16;
defparam dpb_inst_1.BIT_WIDTH_1 = 16;
defparam dpb_inst_1.BLK_SEL_0 = 3'b001;
defparam dpb_inst_1.BLK_SEL_1 = 3'b001;
defparam dpb_inst_1.RESET_MODE = "SYNC";

DPB dpb_inst_2 (
    .DOA(dpb_inst_2_douta[31:16]),
    .DOB(dpb_inst_2_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_2.READ_MODE0 = 1'b0;
defparam dpb_inst_2.READ_MODE1 = 1'b0;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 16;
defparam dpb_inst_2.BIT_WIDTH_1 = 16;
defparam dpb_inst_2.BLK_SEL_0 = 3'b000;
defparam dpb_inst_2.BLK_SEL_1 = 3'b000;
defparam dpb_inst_2.RESET_MODE = "SYNC";

DPB dpb_inst_3 (
    .DOA(dpb_inst_3_douta[31:16]),
    .DOB(dpb_inst_3_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_3.READ_MODE0 = 1'b0;
defparam dpb_inst_3.READ_MODE1 = 1'b0;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 16;
defparam dpb_inst_3.BIT_WIDTH_1 = 16;
defparam dpb_inst_3.BLK_SEL_0 = 3'b001;
defparam dpb_inst_3.BLK_SEL_1 = 3'b001;
defparam dpb_inst_3.RESET_MODE = "SYNC";

DPB dpb_inst_4 (
    .DOA(dpb_inst_4_douta[47:32]),
    .DOB(dpb_inst_4_doutb[47:32]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[47:32]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[47:32])
);

defparam dpb_inst_4.READ_MODE0 = 1'b0;
defparam dpb_inst_4.READ_MODE1 = 1'b0;
defparam dpb_inst_4.WRITE_MODE0 = 2'b00;
defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
defparam dpb_inst_4.BIT_WIDTH_0 = 16;
defparam dpb_inst_4.BIT_WIDTH_1 = 16;
defparam dpb_inst_4.BLK_SEL_0 = 3'b000;
defparam dpb_inst_4.BLK_SEL_1 = 3'b000;
defparam dpb_inst_4.RESET_MODE = "SYNC";

DPB dpb_inst_5 (
    .DOA(dpb_inst_5_douta[47:32]),
    .DOB(dpb_inst_5_doutb[47:32]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[47:32]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[47:32])
);

defparam dpb_inst_5.READ_MODE0 = 1'b0;
defparam dpb_inst_5.READ_MODE1 = 1'b0;
defparam dpb_inst_5.WRITE_MODE0 = 2'b00;
defparam dpb_inst_5.WRITE_MODE1 = 2'b00;
defparam dpb_inst_5.BIT_WIDTH_0 = 16;
defparam dpb_inst_5.BIT_WIDTH_1 = 16;
defparam dpb_inst_5.BLK_SEL_0 = 3'b001;
defparam dpb_inst_5.BLK_SEL_1 = 3'b001;
defparam dpb_inst_5.RESET_MODE = "SYNC";

DPB dpb_inst_6 (
    .DOA(dpb_inst_6_douta[63:48]),
    .DOB(dpb_inst_6_doutb[63:48]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[63:48]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[63:48])
);

defparam dpb_inst_6.READ_MODE0 = 1'b0;
defparam dpb_inst_6.READ_MODE1 = 1'b0;
defparam dpb_inst_6.WRITE_MODE0 = 2'b00;
defparam dpb_inst_6.WRITE_MODE1 = 2'b00;
defparam dpb_inst_6.BIT_WIDTH_0 = 16;
defparam dpb_inst_6.BIT_WIDTH_1 = 16;
defparam dpb_inst_6.BLK_SEL_0 = 3'b000;
defparam dpb_inst_6.BLK_SEL_1 = 3'b000;
defparam dpb_inst_6.RESET_MODE = "SYNC";

DPB dpb_inst_7 (
    .DOA(dpb_inst_7_douta[63:48]),
    .DOB(dpb_inst_7_doutb[63:48]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[63:48]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[63:48])
);

defparam dpb_inst_7.READ_MODE0 = 1'b0;
defparam dpb_inst_7.READ_MODE1 = 1'b0;
defparam dpb_inst_7.WRITE_MODE0 = 2'b00;
defparam dpb_inst_7.WRITE_MODE1 = 2'b00;
defparam dpb_inst_7.BIT_WIDTH_0 = 16;
defparam dpb_inst_7.BIT_WIDTH_1 = 16;
defparam dpb_inst_7.BLK_SEL_0 = 3'b001;
defparam dpb_inst_7.BLK_SEL_1 = 3'b001;
defparam dpb_inst_7.RESET_MODE = "SYNC";

DPB dpb_inst_8 (
    .DOA(dpb_inst_8_douta[79:64]),
    .DOB(dpb_inst_8_doutb[79:64]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[79:64]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[79:64])
);

defparam dpb_inst_8.READ_MODE0 = 1'b0;
defparam dpb_inst_8.READ_MODE1 = 1'b0;
defparam dpb_inst_8.WRITE_MODE0 = 2'b00;
defparam dpb_inst_8.WRITE_MODE1 = 2'b00;
defparam dpb_inst_8.BIT_WIDTH_0 = 16;
defparam dpb_inst_8.BIT_WIDTH_1 = 16;
defparam dpb_inst_8.BLK_SEL_0 = 3'b000;
defparam dpb_inst_8.BLK_SEL_1 = 3'b000;
defparam dpb_inst_8.RESET_MODE = "SYNC";

DPB dpb_inst_9 (
    .DOA(dpb_inst_9_douta[79:64]),
    .DOB(dpb_inst_9_doutb[79:64]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[79:64]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[79:64])
);

defparam dpb_inst_9.READ_MODE0 = 1'b0;
defparam dpb_inst_9.READ_MODE1 = 1'b0;
defparam dpb_inst_9.WRITE_MODE0 = 2'b00;
defparam dpb_inst_9.WRITE_MODE1 = 2'b00;
defparam dpb_inst_9.BIT_WIDTH_0 = 16;
defparam dpb_inst_9.BIT_WIDTH_1 = 16;
defparam dpb_inst_9.BLK_SEL_0 = 3'b001;
defparam dpb_inst_9.BLK_SEL_1 = 3'b001;
defparam dpb_inst_9.RESET_MODE = "SYNC";

DPB dpb_inst_10 (
    .DOA(dpb_inst_10_douta[95:80]),
    .DOB(dpb_inst_10_doutb[95:80]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[95:80]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[95:80])
);

defparam dpb_inst_10.READ_MODE0 = 1'b0;
defparam dpb_inst_10.READ_MODE1 = 1'b0;
defparam dpb_inst_10.WRITE_MODE0 = 2'b00;
defparam dpb_inst_10.WRITE_MODE1 = 2'b00;
defparam dpb_inst_10.BIT_WIDTH_0 = 16;
defparam dpb_inst_10.BIT_WIDTH_1 = 16;
defparam dpb_inst_10.BLK_SEL_0 = 3'b000;
defparam dpb_inst_10.BLK_SEL_1 = 3'b000;
defparam dpb_inst_10.RESET_MODE = "SYNC";

DPB dpb_inst_11 (
    .DOA(dpb_inst_11_douta[95:80]),
    .DOB(dpb_inst_11_doutb[95:80]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[95:80]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[95:80])
);

defparam dpb_inst_11.READ_MODE0 = 1'b0;
defparam dpb_inst_11.READ_MODE1 = 1'b0;
defparam dpb_inst_11.WRITE_MODE0 = 2'b00;
defparam dpb_inst_11.WRITE_MODE1 = 2'b00;
defparam dpb_inst_11.BIT_WIDTH_0 = 16;
defparam dpb_inst_11.BIT_WIDTH_1 = 16;
defparam dpb_inst_11.BLK_SEL_0 = 3'b001;
defparam dpb_inst_11.BLK_SEL_1 = 3'b001;
defparam dpb_inst_11.RESET_MODE = "SYNC";

DPB dpb_inst_12 (
    .DOA(dpb_inst_12_douta[111:96]),
    .DOB(dpb_inst_12_doutb[111:96]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[111:96]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[111:96])
);

defparam dpb_inst_12.READ_MODE0 = 1'b0;
defparam dpb_inst_12.READ_MODE1 = 1'b0;
defparam dpb_inst_12.WRITE_MODE0 = 2'b00;
defparam dpb_inst_12.WRITE_MODE1 = 2'b00;
defparam dpb_inst_12.BIT_WIDTH_0 = 16;
defparam dpb_inst_12.BIT_WIDTH_1 = 16;
defparam dpb_inst_12.BLK_SEL_0 = 3'b000;
defparam dpb_inst_12.BLK_SEL_1 = 3'b000;
defparam dpb_inst_12.RESET_MODE = "SYNC";

DPB dpb_inst_13 (
    .DOA(dpb_inst_13_douta[111:96]),
    .DOB(dpb_inst_13_doutb[111:96]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[111:96]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[111:96])
);

defparam dpb_inst_13.READ_MODE0 = 1'b0;
defparam dpb_inst_13.READ_MODE1 = 1'b0;
defparam dpb_inst_13.WRITE_MODE0 = 2'b00;
defparam dpb_inst_13.WRITE_MODE1 = 2'b00;
defparam dpb_inst_13.BIT_WIDTH_0 = 16;
defparam dpb_inst_13.BIT_WIDTH_1 = 16;
defparam dpb_inst_13.BLK_SEL_0 = 3'b001;
defparam dpb_inst_13.BLK_SEL_1 = 3'b001;
defparam dpb_inst_13.RESET_MODE = "SYNC";

DPB dpb_inst_14 (
    .DOA(dpb_inst_14_douta[127:112]),
    .DOB(dpb_inst_14_doutb[127:112]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[127:112]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[127:112])
);

defparam dpb_inst_14.READ_MODE0 = 1'b0;
defparam dpb_inst_14.READ_MODE1 = 1'b0;
defparam dpb_inst_14.WRITE_MODE0 = 2'b00;
defparam dpb_inst_14.WRITE_MODE1 = 2'b00;
defparam dpb_inst_14.BIT_WIDTH_0 = 16;
defparam dpb_inst_14.BIT_WIDTH_1 = 16;
defparam dpb_inst_14.BLK_SEL_0 = 3'b000;
defparam dpb_inst_14.BLK_SEL_1 = 3'b000;
defparam dpb_inst_14.RESET_MODE = "SYNC";

DPB dpb_inst_15 (
    .DOA(dpb_inst_15_douta[127:112]),
    .DOB(dpb_inst_15_doutb[127:112]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[10]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIA(dina[127:112]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DIB(dinb[127:112])
);

defparam dpb_inst_15.READ_MODE0 = 1'b0;
defparam dpb_inst_15.READ_MODE1 = 1'b0;
defparam dpb_inst_15.WRITE_MODE0 = 2'b00;
defparam dpb_inst_15.WRITE_MODE1 = 2'b00;
defparam dpb_inst_15.BIT_WIDTH_0 = 16;
defparam dpb_inst_15.BIT_WIDTH_1 = 16;
defparam dpb_inst_15.BLK_SEL_0 = 3'b001;
defparam dpb_inst_15.BLK_SEL_1 = 3'b001;
defparam dpb_inst_15.RESET_MODE = "SYNC";

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[10]),
  .CLK(clka),
  .CE(cea_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[10]),
  .CLK(clkb),
  .CE(ceb_w)
);
MUX2 mux_inst_0 (
  .O(douta[0]),
  .I0(dpb_inst_0_douta[0]),
  .I1(dpb_inst_1_douta[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_1 (
  .O(douta[1]),
  .I0(dpb_inst_0_douta[1]),
  .I1(dpb_inst_1_douta[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_2 (
  .O(douta[2]),
  .I0(dpb_inst_0_douta[2]),
  .I1(dpb_inst_1_douta[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_3 (
  .O(douta[3]),
  .I0(dpb_inst_0_douta[3]),
  .I1(dpb_inst_1_douta[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_4 (
  .O(douta[4]),
  .I0(dpb_inst_0_douta[4]),
  .I1(dpb_inst_1_douta[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(douta[5]),
  .I0(dpb_inst_0_douta[5]),
  .I1(dpb_inst_1_douta[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_6 (
  .O(douta[6]),
  .I0(dpb_inst_0_douta[6]),
  .I1(dpb_inst_1_douta[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_7 (
  .O(douta[7]),
  .I0(dpb_inst_0_douta[7]),
  .I1(dpb_inst_1_douta[7]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(douta[8]),
  .I0(dpb_inst_0_douta[8]),
  .I1(dpb_inst_1_douta[8]),
  .S0(dff_q_0)
);
MUX2 mux_inst_9 (
  .O(douta[9]),
  .I0(dpb_inst_0_douta[9]),
  .I1(dpb_inst_1_douta[9]),
  .S0(dff_q_0)
);
MUX2 mux_inst_10 (
  .O(douta[10]),
  .I0(dpb_inst_0_douta[10]),
  .I1(dpb_inst_1_douta[10]),
  .S0(dff_q_0)
);
MUX2 mux_inst_11 (
  .O(douta[11]),
  .I0(dpb_inst_0_douta[11]),
  .I1(dpb_inst_1_douta[11]),
  .S0(dff_q_0)
);
MUX2 mux_inst_12 (
  .O(douta[12]),
  .I0(dpb_inst_0_douta[12]),
  .I1(dpb_inst_1_douta[12]),
  .S0(dff_q_0)
);
MUX2 mux_inst_13 (
  .O(douta[13]),
  .I0(dpb_inst_0_douta[13]),
  .I1(dpb_inst_1_douta[13]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(douta[14]),
  .I0(dpb_inst_0_douta[14]),
  .I1(dpb_inst_1_douta[14]),
  .S0(dff_q_0)
);
MUX2 mux_inst_15 (
  .O(douta[15]),
  .I0(dpb_inst_0_douta[15]),
  .I1(dpb_inst_1_douta[15]),
  .S0(dff_q_0)
);
MUX2 mux_inst_16 (
  .O(douta[16]),
  .I0(dpb_inst_2_douta[16]),
  .I1(dpb_inst_3_douta[16]),
  .S0(dff_q_0)
);
MUX2 mux_inst_17 (
  .O(douta[17]),
  .I0(dpb_inst_2_douta[17]),
  .I1(dpb_inst_3_douta[17]),
  .S0(dff_q_0)
);
MUX2 mux_inst_18 (
  .O(douta[18]),
  .I0(dpb_inst_2_douta[18]),
  .I1(dpb_inst_3_douta[18]),
  .S0(dff_q_0)
);
MUX2 mux_inst_19 (
  .O(douta[19]),
  .I0(dpb_inst_2_douta[19]),
  .I1(dpb_inst_3_douta[19]),
  .S0(dff_q_0)
);
MUX2 mux_inst_20 (
  .O(douta[20]),
  .I0(dpb_inst_2_douta[20]),
  .I1(dpb_inst_3_douta[20]),
  .S0(dff_q_0)
);
MUX2 mux_inst_21 (
  .O(douta[21]),
  .I0(dpb_inst_2_douta[21]),
  .I1(dpb_inst_3_douta[21]),
  .S0(dff_q_0)
);
MUX2 mux_inst_22 (
  .O(douta[22]),
  .I0(dpb_inst_2_douta[22]),
  .I1(dpb_inst_3_douta[22]),
  .S0(dff_q_0)
);
MUX2 mux_inst_23 (
  .O(douta[23]),
  .I0(dpb_inst_2_douta[23]),
  .I1(dpb_inst_3_douta[23]),
  .S0(dff_q_0)
);
MUX2 mux_inst_24 (
  .O(douta[24]),
  .I0(dpb_inst_2_douta[24]),
  .I1(dpb_inst_3_douta[24]),
  .S0(dff_q_0)
);
MUX2 mux_inst_25 (
  .O(douta[25]),
  .I0(dpb_inst_2_douta[25]),
  .I1(dpb_inst_3_douta[25]),
  .S0(dff_q_0)
);
MUX2 mux_inst_26 (
  .O(douta[26]),
  .I0(dpb_inst_2_douta[26]),
  .I1(dpb_inst_3_douta[26]),
  .S0(dff_q_0)
);
MUX2 mux_inst_27 (
  .O(douta[27]),
  .I0(dpb_inst_2_douta[27]),
  .I1(dpb_inst_3_douta[27]),
  .S0(dff_q_0)
);
MUX2 mux_inst_28 (
  .O(douta[28]),
  .I0(dpb_inst_2_douta[28]),
  .I1(dpb_inst_3_douta[28]),
  .S0(dff_q_0)
);
MUX2 mux_inst_29 (
  .O(douta[29]),
  .I0(dpb_inst_2_douta[29]),
  .I1(dpb_inst_3_douta[29]),
  .S0(dff_q_0)
);
MUX2 mux_inst_30 (
  .O(douta[30]),
  .I0(dpb_inst_2_douta[30]),
  .I1(dpb_inst_3_douta[30]),
  .S0(dff_q_0)
);
MUX2 mux_inst_31 (
  .O(douta[31]),
  .I0(dpb_inst_2_douta[31]),
  .I1(dpb_inst_3_douta[31]),
  .S0(dff_q_0)
);
MUX2 mux_inst_32 (
  .O(douta[32]),
  .I0(dpb_inst_4_douta[32]),
  .I1(dpb_inst_5_douta[32]),
  .S0(dff_q_0)
);
MUX2 mux_inst_33 (
  .O(douta[33]),
  .I0(dpb_inst_4_douta[33]),
  .I1(dpb_inst_5_douta[33]),
  .S0(dff_q_0)
);
MUX2 mux_inst_34 (
  .O(douta[34]),
  .I0(dpb_inst_4_douta[34]),
  .I1(dpb_inst_5_douta[34]),
  .S0(dff_q_0)
);
MUX2 mux_inst_35 (
  .O(douta[35]),
  .I0(dpb_inst_4_douta[35]),
  .I1(dpb_inst_5_douta[35]),
  .S0(dff_q_0)
);
MUX2 mux_inst_36 (
  .O(douta[36]),
  .I0(dpb_inst_4_douta[36]),
  .I1(dpb_inst_5_douta[36]),
  .S0(dff_q_0)
);
MUX2 mux_inst_37 (
  .O(douta[37]),
  .I0(dpb_inst_4_douta[37]),
  .I1(dpb_inst_5_douta[37]),
  .S0(dff_q_0)
);
MUX2 mux_inst_38 (
  .O(douta[38]),
  .I0(dpb_inst_4_douta[38]),
  .I1(dpb_inst_5_douta[38]),
  .S0(dff_q_0)
);
MUX2 mux_inst_39 (
  .O(douta[39]),
  .I0(dpb_inst_4_douta[39]),
  .I1(dpb_inst_5_douta[39]),
  .S0(dff_q_0)
);
MUX2 mux_inst_40 (
  .O(douta[40]),
  .I0(dpb_inst_4_douta[40]),
  .I1(dpb_inst_5_douta[40]),
  .S0(dff_q_0)
);
MUX2 mux_inst_41 (
  .O(douta[41]),
  .I0(dpb_inst_4_douta[41]),
  .I1(dpb_inst_5_douta[41]),
  .S0(dff_q_0)
);
MUX2 mux_inst_42 (
  .O(douta[42]),
  .I0(dpb_inst_4_douta[42]),
  .I1(dpb_inst_5_douta[42]),
  .S0(dff_q_0)
);
MUX2 mux_inst_43 (
  .O(douta[43]),
  .I0(dpb_inst_4_douta[43]),
  .I1(dpb_inst_5_douta[43]),
  .S0(dff_q_0)
);
MUX2 mux_inst_44 (
  .O(douta[44]),
  .I0(dpb_inst_4_douta[44]),
  .I1(dpb_inst_5_douta[44]),
  .S0(dff_q_0)
);
MUX2 mux_inst_45 (
  .O(douta[45]),
  .I0(dpb_inst_4_douta[45]),
  .I1(dpb_inst_5_douta[45]),
  .S0(dff_q_0)
);
MUX2 mux_inst_46 (
  .O(douta[46]),
  .I0(dpb_inst_4_douta[46]),
  .I1(dpb_inst_5_douta[46]),
  .S0(dff_q_0)
);
MUX2 mux_inst_47 (
  .O(douta[47]),
  .I0(dpb_inst_4_douta[47]),
  .I1(dpb_inst_5_douta[47]),
  .S0(dff_q_0)
);
MUX2 mux_inst_48 (
  .O(douta[48]),
  .I0(dpb_inst_6_douta[48]),
  .I1(dpb_inst_7_douta[48]),
  .S0(dff_q_0)
);
MUX2 mux_inst_49 (
  .O(douta[49]),
  .I0(dpb_inst_6_douta[49]),
  .I1(dpb_inst_7_douta[49]),
  .S0(dff_q_0)
);
MUX2 mux_inst_50 (
  .O(douta[50]),
  .I0(dpb_inst_6_douta[50]),
  .I1(dpb_inst_7_douta[50]),
  .S0(dff_q_0)
);
MUX2 mux_inst_51 (
  .O(douta[51]),
  .I0(dpb_inst_6_douta[51]),
  .I1(dpb_inst_7_douta[51]),
  .S0(dff_q_0)
);
MUX2 mux_inst_52 (
  .O(douta[52]),
  .I0(dpb_inst_6_douta[52]),
  .I1(dpb_inst_7_douta[52]),
  .S0(dff_q_0)
);
MUX2 mux_inst_53 (
  .O(douta[53]),
  .I0(dpb_inst_6_douta[53]),
  .I1(dpb_inst_7_douta[53]),
  .S0(dff_q_0)
);
MUX2 mux_inst_54 (
  .O(douta[54]),
  .I0(dpb_inst_6_douta[54]),
  .I1(dpb_inst_7_douta[54]),
  .S0(dff_q_0)
);
MUX2 mux_inst_55 (
  .O(douta[55]),
  .I0(dpb_inst_6_douta[55]),
  .I1(dpb_inst_7_douta[55]),
  .S0(dff_q_0)
);
MUX2 mux_inst_56 (
  .O(douta[56]),
  .I0(dpb_inst_6_douta[56]),
  .I1(dpb_inst_7_douta[56]),
  .S0(dff_q_0)
);
MUX2 mux_inst_57 (
  .O(douta[57]),
  .I0(dpb_inst_6_douta[57]),
  .I1(dpb_inst_7_douta[57]),
  .S0(dff_q_0)
);
MUX2 mux_inst_58 (
  .O(douta[58]),
  .I0(dpb_inst_6_douta[58]),
  .I1(dpb_inst_7_douta[58]),
  .S0(dff_q_0)
);
MUX2 mux_inst_59 (
  .O(douta[59]),
  .I0(dpb_inst_6_douta[59]),
  .I1(dpb_inst_7_douta[59]),
  .S0(dff_q_0)
);
MUX2 mux_inst_60 (
  .O(douta[60]),
  .I0(dpb_inst_6_douta[60]),
  .I1(dpb_inst_7_douta[60]),
  .S0(dff_q_0)
);
MUX2 mux_inst_61 (
  .O(douta[61]),
  .I0(dpb_inst_6_douta[61]),
  .I1(dpb_inst_7_douta[61]),
  .S0(dff_q_0)
);
MUX2 mux_inst_62 (
  .O(douta[62]),
  .I0(dpb_inst_6_douta[62]),
  .I1(dpb_inst_7_douta[62]),
  .S0(dff_q_0)
);
MUX2 mux_inst_63 (
  .O(douta[63]),
  .I0(dpb_inst_6_douta[63]),
  .I1(dpb_inst_7_douta[63]),
  .S0(dff_q_0)
);
MUX2 mux_inst_64 (
  .O(douta[64]),
  .I0(dpb_inst_8_douta[64]),
  .I1(dpb_inst_9_douta[64]),
  .S0(dff_q_0)
);
MUX2 mux_inst_65 (
  .O(douta[65]),
  .I0(dpb_inst_8_douta[65]),
  .I1(dpb_inst_9_douta[65]),
  .S0(dff_q_0)
);
MUX2 mux_inst_66 (
  .O(douta[66]),
  .I0(dpb_inst_8_douta[66]),
  .I1(dpb_inst_9_douta[66]),
  .S0(dff_q_0)
);
MUX2 mux_inst_67 (
  .O(douta[67]),
  .I0(dpb_inst_8_douta[67]),
  .I1(dpb_inst_9_douta[67]),
  .S0(dff_q_0)
);
MUX2 mux_inst_68 (
  .O(douta[68]),
  .I0(dpb_inst_8_douta[68]),
  .I1(dpb_inst_9_douta[68]),
  .S0(dff_q_0)
);
MUX2 mux_inst_69 (
  .O(douta[69]),
  .I0(dpb_inst_8_douta[69]),
  .I1(dpb_inst_9_douta[69]),
  .S0(dff_q_0)
);
MUX2 mux_inst_70 (
  .O(douta[70]),
  .I0(dpb_inst_8_douta[70]),
  .I1(dpb_inst_9_douta[70]),
  .S0(dff_q_0)
);
MUX2 mux_inst_71 (
  .O(douta[71]),
  .I0(dpb_inst_8_douta[71]),
  .I1(dpb_inst_9_douta[71]),
  .S0(dff_q_0)
);
MUX2 mux_inst_72 (
  .O(douta[72]),
  .I0(dpb_inst_8_douta[72]),
  .I1(dpb_inst_9_douta[72]),
  .S0(dff_q_0)
);
MUX2 mux_inst_73 (
  .O(douta[73]),
  .I0(dpb_inst_8_douta[73]),
  .I1(dpb_inst_9_douta[73]),
  .S0(dff_q_0)
);
MUX2 mux_inst_74 (
  .O(douta[74]),
  .I0(dpb_inst_8_douta[74]),
  .I1(dpb_inst_9_douta[74]),
  .S0(dff_q_0)
);
MUX2 mux_inst_75 (
  .O(douta[75]),
  .I0(dpb_inst_8_douta[75]),
  .I1(dpb_inst_9_douta[75]),
  .S0(dff_q_0)
);
MUX2 mux_inst_76 (
  .O(douta[76]),
  .I0(dpb_inst_8_douta[76]),
  .I1(dpb_inst_9_douta[76]),
  .S0(dff_q_0)
);
MUX2 mux_inst_77 (
  .O(douta[77]),
  .I0(dpb_inst_8_douta[77]),
  .I1(dpb_inst_9_douta[77]),
  .S0(dff_q_0)
);
MUX2 mux_inst_78 (
  .O(douta[78]),
  .I0(dpb_inst_8_douta[78]),
  .I1(dpb_inst_9_douta[78]),
  .S0(dff_q_0)
);
MUX2 mux_inst_79 (
  .O(douta[79]),
  .I0(dpb_inst_8_douta[79]),
  .I1(dpb_inst_9_douta[79]),
  .S0(dff_q_0)
);
MUX2 mux_inst_80 (
  .O(douta[80]),
  .I0(dpb_inst_10_douta[80]),
  .I1(dpb_inst_11_douta[80]),
  .S0(dff_q_0)
);
MUX2 mux_inst_81 (
  .O(douta[81]),
  .I0(dpb_inst_10_douta[81]),
  .I1(dpb_inst_11_douta[81]),
  .S0(dff_q_0)
);
MUX2 mux_inst_82 (
  .O(douta[82]),
  .I0(dpb_inst_10_douta[82]),
  .I1(dpb_inst_11_douta[82]),
  .S0(dff_q_0)
);
MUX2 mux_inst_83 (
  .O(douta[83]),
  .I0(dpb_inst_10_douta[83]),
  .I1(dpb_inst_11_douta[83]),
  .S0(dff_q_0)
);
MUX2 mux_inst_84 (
  .O(douta[84]),
  .I0(dpb_inst_10_douta[84]),
  .I1(dpb_inst_11_douta[84]),
  .S0(dff_q_0)
);
MUX2 mux_inst_85 (
  .O(douta[85]),
  .I0(dpb_inst_10_douta[85]),
  .I1(dpb_inst_11_douta[85]),
  .S0(dff_q_0)
);
MUX2 mux_inst_86 (
  .O(douta[86]),
  .I0(dpb_inst_10_douta[86]),
  .I1(dpb_inst_11_douta[86]),
  .S0(dff_q_0)
);
MUX2 mux_inst_87 (
  .O(douta[87]),
  .I0(dpb_inst_10_douta[87]),
  .I1(dpb_inst_11_douta[87]),
  .S0(dff_q_0)
);
MUX2 mux_inst_88 (
  .O(douta[88]),
  .I0(dpb_inst_10_douta[88]),
  .I1(dpb_inst_11_douta[88]),
  .S0(dff_q_0)
);
MUX2 mux_inst_89 (
  .O(douta[89]),
  .I0(dpb_inst_10_douta[89]),
  .I1(dpb_inst_11_douta[89]),
  .S0(dff_q_0)
);
MUX2 mux_inst_90 (
  .O(douta[90]),
  .I0(dpb_inst_10_douta[90]),
  .I1(dpb_inst_11_douta[90]),
  .S0(dff_q_0)
);
MUX2 mux_inst_91 (
  .O(douta[91]),
  .I0(dpb_inst_10_douta[91]),
  .I1(dpb_inst_11_douta[91]),
  .S0(dff_q_0)
);
MUX2 mux_inst_92 (
  .O(douta[92]),
  .I0(dpb_inst_10_douta[92]),
  .I1(dpb_inst_11_douta[92]),
  .S0(dff_q_0)
);
MUX2 mux_inst_93 (
  .O(douta[93]),
  .I0(dpb_inst_10_douta[93]),
  .I1(dpb_inst_11_douta[93]),
  .S0(dff_q_0)
);
MUX2 mux_inst_94 (
  .O(douta[94]),
  .I0(dpb_inst_10_douta[94]),
  .I1(dpb_inst_11_douta[94]),
  .S0(dff_q_0)
);
MUX2 mux_inst_95 (
  .O(douta[95]),
  .I0(dpb_inst_10_douta[95]),
  .I1(dpb_inst_11_douta[95]),
  .S0(dff_q_0)
);
MUX2 mux_inst_96 (
  .O(douta[96]),
  .I0(dpb_inst_12_douta[96]),
  .I1(dpb_inst_13_douta[96]),
  .S0(dff_q_0)
);
MUX2 mux_inst_97 (
  .O(douta[97]),
  .I0(dpb_inst_12_douta[97]),
  .I1(dpb_inst_13_douta[97]),
  .S0(dff_q_0)
);
MUX2 mux_inst_98 (
  .O(douta[98]),
  .I0(dpb_inst_12_douta[98]),
  .I1(dpb_inst_13_douta[98]),
  .S0(dff_q_0)
);
MUX2 mux_inst_99 (
  .O(douta[99]),
  .I0(dpb_inst_12_douta[99]),
  .I1(dpb_inst_13_douta[99]),
  .S0(dff_q_0)
);
MUX2 mux_inst_100 (
  .O(douta[100]),
  .I0(dpb_inst_12_douta[100]),
  .I1(dpb_inst_13_douta[100]),
  .S0(dff_q_0)
);
MUX2 mux_inst_101 (
  .O(douta[101]),
  .I0(dpb_inst_12_douta[101]),
  .I1(dpb_inst_13_douta[101]),
  .S0(dff_q_0)
);
MUX2 mux_inst_102 (
  .O(douta[102]),
  .I0(dpb_inst_12_douta[102]),
  .I1(dpb_inst_13_douta[102]),
  .S0(dff_q_0)
);
MUX2 mux_inst_103 (
  .O(douta[103]),
  .I0(dpb_inst_12_douta[103]),
  .I1(dpb_inst_13_douta[103]),
  .S0(dff_q_0)
);
MUX2 mux_inst_104 (
  .O(douta[104]),
  .I0(dpb_inst_12_douta[104]),
  .I1(dpb_inst_13_douta[104]),
  .S0(dff_q_0)
);
MUX2 mux_inst_105 (
  .O(douta[105]),
  .I0(dpb_inst_12_douta[105]),
  .I1(dpb_inst_13_douta[105]),
  .S0(dff_q_0)
);
MUX2 mux_inst_106 (
  .O(douta[106]),
  .I0(dpb_inst_12_douta[106]),
  .I1(dpb_inst_13_douta[106]),
  .S0(dff_q_0)
);
MUX2 mux_inst_107 (
  .O(douta[107]),
  .I0(dpb_inst_12_douta[107]),
  .I1(dpb_inst_13_douta[107]),
  .S0(dff_q_0)
);
MUX2 mux_inst_108 (
  .O(douta[108]),
  .I0(dpb_inst_12_douta[108]),
  .I1(dpb_inst_13_douta[108]),
  .S0(dff_q_0)
);
MUX2 mux_inst_109 (
  .O(douta[109]),
  .I0(dpb_inst_12_douta[109]),
  .I1(dpb_inst_13_douta[109]),
  .S0(dff_q_0)
);
MUX2 mux_inst_110 (
  .O(douta[110]),
  .I0(dpb_inst_12_douta[110]),
  .I1(dpb_inst_13_douta[110]),
  .S0(dff_q_0)
);
MUX2 mux_inst_111 (
  .O(douta[111]),
  .I0(dpb_inst_12_douta[111]),
  .I1(dpb_inst_13_douta[111]),
  .S0(dff_q_0)
);
MUX2 mux_inst_112 (
  .O(douta[112]),
  .I0(dpb_inst_14_douta[112]),
  .I1(dpb_inst_15_douta[112]),
  .S0(dff_q_0)
);
MUX2 mux_inst_113 (
  .O(douta[113]),
  .I0(dpb_inst_14_douta[113]),
  .I1(dpb_inst_15_douta[113]),
  .S0(dff_q_0)
);
MUX2 mux_inst_114 (
  .O(douta[114]),
  .I0(dpb_inst_14_douta[114]),
  .I1(dpb_inst_15_douta[114]),
  .S0(dff_q_0)
);
MUX2 mux_inst_115 (
  .O(douta[115]),
  .I0(dpb_inst_14_douta[115]),
  .I1(dpb_inst_15_douta[115]),
  .S0(dff_q_0)
);
MUX2 mux_inst_116 (
  .O(douta[116]),
  .I0(dpb_inst_14_douta[116]),
  .I1(dpb_inst_15_douta[116]),
  .S0(dff_q_0)
);
MUX2 mux_inst_117 (
  .O(douta[117]),
  .I0(dpb_inst_14_douta[117]),
  .I1(dpb_inst_15_douta[117]),
  .S0(dff_q_0)
);
MUX2 mux_inst_118 (
  .O(douta[118]),
  .I0(dpb_inst_14_douta[118]),
  .I1(dpb_inst_15_douta[118]),
  .S0(dff_q_0)
);
MUX2 mux_inst_119 (
  .O(douta[119]),
  .I0(dpb_inst_14_douta[119]),
  .I1(dpb_inst_15_douta[119]),
  .S0(dff_q_0)
);
MUX2 mux_inst_120 (
  .O(douta[120]),
  .I0(dpb_inst_14_douta[120]),
  .I1(dpb_inst_15_douta[120]),
  .S0(dff_q_0)
);
MUX2 mux_inst_121 (
  .O(douta[121]),
  .I0(dpb_inst_14_douta[121]),
  .I1(dpb_inst_15_douta[121]),
  .S0(dff_q_0)
);
MUX2 mux_inst_122 (
  .O(douta[122]),
  .I0(dpb_inst_14_douta[122]),
  .I1(dpb_inst_15_douta[122]),
  .S0(dff_q_0)
);
MUX2 mux_inst_123 (
  .O(douta[123]),
  .I0(dpb_inst_14_douta[123]),
  .I1(dpb_inst_15_douta[123]),
  .S0(dff_q_0)
);
MUX2 mux_inst_124 (
  .O(douta[124]),
  .I0(dpb_inst_14_douta[124]),
  .I1(dpb_inst_15_douta[124]),
  .S0(dff_q_0)
);
MUX2 mux_inst_125 (
  .O(douta[125]),
  .I0(dpb_inst_14_douta[125]),
  .I1(dpb_inst_15_douta[125]),
  .S0(dff_q_0)
);
MUX2 mux_inst_126 (
  .O(douta[126]),
  .I0(dpb_inst_14_douta[126]),
  .I1(dpb_inst_15_douta[126]),
  .S0(dff_q_0)
);
MUX2 mux_inst_127 (
  .O(douta[127]),
  .I0(dpb_inst_14_douta[127]),
  .I1(dpb_inst_15_douta[127]),
  .S0(dff_q_0)
);
MUX2 mux_inst_128 (
  .O(doutb[0]),
  .I0(dpb_inst_0_doutb[0]),
  .I1(dpb_inst_1_doutb[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_129 (
  .O(doutb[1]),
  .I0(dpb_inst_0_doutb[1]),
  .I1(dpb_inst_1_doutb[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_130 (
  .O(doutb[2]),
  .I0(dpb_inst_0_doutb[2]),
  .I1(dpb_inst_1_doutb[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_131 (
  .O(doutb[3]),
  .I0(dpb_inst_0_doutb[3]),
  .I1(dpb_inst_1_doutb[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_132 (
  .O(doutb[4]),
  .I0(dpb_inst_0_doutb[4]),
  .I1(dpb_inst_1_doutb[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_133 (
  .O(doutb[5]),
  .I0(dpb_inst_0_doutb[5]),
  .I1(dpb_inst_1_doutb[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_134 (
  .O(doutb[6]),
  .I0(dpb_inst_0_doutb[6]),
  .I1(dpb_inst_1_doutb[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_135 (
  .O(doutb[7]),
  .I0(dpb_inst_0_doutb[7]),
  .I1(dpb_inst_1_doutb[7]),
  .S0(dff_q_1)
);
MUX2 mux_inst_136 (
  .O(doutb[8]),
  .I0(dpb_inst_0_doutb[8]),
  .I1(dpb_inst_1_doutb[8]),
  .S0(dff_q_1)
);
MUX2 mux_inst_137 (
  .O(doutb[9]),
  .I0(dpb_inst_0_doutb[9]),
  .I1(dpb_inst_1_doutb[9]),
  .S0(dff_q_1)
);
MUX2 mux_inst_138 (
  .O(doutb[10]),
  .I0(dpb_inst_0_doutb[10]),
  .I1(dpb_inst_1_doutb[10]),
  .S0(dff_q_1)
);
MUX2 mux_inst_139 (
  .O(doutb[11]),
  .I0(dpb_inst_0_doutb[11]),
  .I1(dpb_inst_1_doutb[11]),
  .S0(dff_q_1)
);
MUX2 mux_inst_140 (
  .O(doutb[12]),
  .I0(dpb_inst_0_doutb[12]),
  .I1(dpb_inst_1_doutb[12]),
  .S0(dff_q_1)
);
MUX2 mux_inst_141 (
  .O(doutb[13]),
  .I0(dpb_inst_0_doutb[13]),
  .I1(dpb_inst_1_doutb[13]),
  .S0(dff_q_1)
);
MUX2 mux_inst_142 (
  .O(doutb[14]),
  .I0(dpb_inst_0_doutb[14]),
  .I1(dpb_inst_1_doutb[14]),
  .S0(dff_q_1)
);
MUX2 mux_inst_143 (
  .O(doutb[15]),
  .I0(dpb_inst_0_doutb[15]),
  .I1(dpb_inst_1_doutb[15]),
  .S0(dff_q_1)
);
MUX2 mux_inst_144 (
  .O(doutb[16]),
  .I0(dpb_inst_2_doutb[16]),
  .I1(dpb_inst_3_doutb[16]),
  .S0(dff_q_1)
);
MUX2 mux_inst_145 (
  .O(doutb[17]),
  .I0(dpb_inst_2_doutb[17]),
  .I1(dpb_inst_3_doutb[17]),
  .S0(dff_q_1)
);
MUX2 mux_inst_146 (
  .O(doutb[18]),
  .I0(dpb_inst_2_doutb[18]),
  .I1(dpb_inst_3_doutb[18]),
  .S0(dff_q_1)
);
MUX2 mux_inst_147 (
  .O(doutb[19]),
  .I0(dpb_inst_2_doutb[19]),
  .I1(dpb_inst_3_doutb[19]),
  .S0(dff_q_1)
);
MUX2 mux_inst_148 (
  .O(doutb[20]),
  .I0(dpb_inst_2_doutb[20]),
  .I1(dpb_inst_3_doutb[20]),
  .S0(dff_q_1)
);
MUX2 mux_inst_149 (
  .O(doutb[21]),
  .I0(dpb_inst_2_doutb[21]),
  .I1(dpb_inst_3_doutb[21]),
  .S0(dff_q_1)
);
MUX2 mux_inst_150 (
  .O(doutb[22]),
  .I0(dpb_inst_2_doutb[22]),
  .I1(dpb_inst_3_doutb[22]),
  .S0(dff_q_1)
);
MUX2 mux_inst_151 (
  .O(doutb[23]),
  .I0(dpb_inst_2_doutb[23]),
  .I1(dpb_inst_3_doutb[23]),
  .S0(dff_q_1)
);
MUX2 mux_inst_152 (
  .O(doutb[24]),
  .I0(dpb_inst_2_doutb[24]),
  .I1(dpb_inst_3_doutb[24]),
  .S0(dff_q_1)
);
MUX2 mux_inst_153 (
  .O(doutb[25]),
  .I0(dpb_inst_2_doutb[25]),
  .I1(dpb_inst_3_doutb[25]),
  .S0(dff_q_1)
);
MUX2 mux_inst_154 (
  .O(doutb[26]),
  .I0(dpb_inst_2_doutb[26]),
  .I1(dpb_inst_3_doutb[26]),
  .S0(dff_q_1)
);
MUX2 mux_inst_155 (
  .O(doutb[27]),
  .I0(dpb_inst_2_doutb[27]),
  .I1(dpb_inst_3_doutb[27]),
  .S0(dff_q_1)
);
MUX2 mux_inst_156 (
  .O(doutb[28]),
  .I0(dpb_inst_2_doutb[28]),
  .I1(dpb_inst_3_doutb[28]),
  .S0(dff_q_1)
);
MUX2 mux_inst_157 (
  .O(doutb[29]),
  .I0(dpb_inst_2_doutb[29]),
  .I1(dpb_inst_3_doutb[29]),
  .S0(dff_q_1)
);
MUX2 mux_inst_158 (
  .O(doutb[30]),
  .I0(dpb_inst_2_doutb[30]),
  .I1(dpb_inst_3_doutb[30]),
  .S0(dff_q_1)
);
MUX2 mux_inst_159 (
  .O(doutb[31]),
  .I0(dpb_inst_2_doutb[31]),
  .I1(dpb_inst_3_doutb[31]),
  .S0(dff_q_1)
);
MUX2 mux_inst_160 (
  .O(doutb[32]),
  .I0(dpb_inst_4_doutb[32]),
  .I1(dpb_inst_5_doutb[32]),
  .S0(dff_q_1)
);
MUX2 mux_inst_161 (
  .O(doutb[33]),
  .I0(dpb_inst_4_doutb[33]),
  .I1(dpb_inst_5_doutb[33]),
  .S0(dff_q_1)
);
MUX2 mux_inst_162 (
  .O(doutb[34]),
  .I0(dpb_inst_4_doutb[34]),
  .I1(dpb_inst_5_doutb[34]),
  .S0(dff_q_1)
);
MUX2 mux_inst_163 (
  .O(doutb[35]),
  .I0(dpb_inst_4_doutb[35]),
  .I1(dpb_inst_5_doutb[35]),
  .S0(dff_q_1)
);
MUX2 mux_inst_164 (
  .O(doutb[36]),
  .I0(dpb_inst_4_doutb[36]),
  .I1(dpb_inst_5_doutb[36]),
  .S0(dff_q_1)
);
MUX2 mux_inst_165 (
  .O(doutb[37]),
  .I0(dpb_inst_4_doutb[37]),
  .I1(dpb_inst_5_doutb[37]),
  .S0(dff_q_1)
);
MUX2 mux_inst_166 (
  .O(doutb[38]),
  .I0(dpb_inst_4_doutb[38]),
  .I1(dpb_inst_5_doutb[38]),
  .S0(dff_q_1)
);
MUX2 mux_inst_167 (
  .O(doutb[39]),
  .I0(dpb_inst_4_doutb[39]),
  .I1(dpb_inst_5_doutb[39]),
  .S0(dff_q_1)
);
MUX2 mux_inst_168 (
  .O(doutb[40]),
  .I0(dpb_inst_4_doutb[40]),
  .I1(dpb_inst_5_doutb[40]),
  .S0(dff_q_1)
);
MUX2 mux_inst_169 (
  .O(doutb[41]),
  .I0(dpb_inst_4_doutb[41]),
  .I1(dpb_inst_5_doutb[41]),
  .S0(dff_q_1)
);
MUX2 mux_inst_170 (
  .O(doutb[42]),
  .I0(dpb_inst_4_doutb[42]),
  .I1(dpb_inst_5_doutb[42]),
  .S0(dff_q_1)
);
MUX2 mux_inst_171 (
  .O(doutb[43]),
  .I0(dpb_inst_4_doutb[43]),
  .I1(dpb_inst_5_doutb[43]),
  .S0(dff_q_1)
);
MUX2 mux_inst_172 (
  .O(doutb[44]),
  .I0(dpb_inst_4_doutb[44]),
  .I1(dpb_inst_5_doutb[44]),
  .S0(dff_q_1)
);
MUX2 mux_inst_173 (
  .O(doutb[45]),
  .I0(dpb_inst_4_doutb[45]),
  .I1(dpb_inst_5_doutb[45]),
  .S0(dff_q_1)
);
MUX2 mux_inst_174 (
  .O(doutb[46]),
  .I0(dpb_inst_4_doutb[46]),
  .I1(dpb_inst_5_doutb[46]),
  .S0(dff_q_1)
);
MUX2 mux_inst_175 (
  .O(doutb[47]),
  .I0(dpb_inst_4_doutb[47]),
  .I1(dpb_inst_5_doutb[47]),
  .S0(dff_q_1)
);
MUX2 mux_inst_176 (
  .O(doutb[48]),
  .I0(dpb_inst_6_doutb[48]),
  .I1(dpb_inst_7_doutb[48]),
  .S0(dff_q_1)
);
MUX2 mux_inst_177 (
  .O(doutb[49]),
  .I0(dpb_inst_6_doutb[49]),
  .I1(dpb_inst_7_doutb[49]),
  .S0(dff_q_1)
);
MUX2 mux_inst_178 (
  .O(doutb[50]),
  .I0(dpb_inst_6_doutb[50]),
  .I1(dpb_inst_7_doutb[50]),
  .S0(dff_q_1)
);
MUX2 mux_inst_179 (
  .O(doutb[51]),
  .I0(dpb_inst_6_doutb[51]),
  .I1(dpb_inst_7_doutb[51]),
  .S0(dff_q_1)
);
MUX2 mux_inst_180 (
  .O(doutb[52]),
  .I0(dpb_inst_6_doutb[52]),
  .I1(dpb_inst_7_doutb[52]),
  .S0(dff_q_1)
);
MUX2 mux_inst_181 (
  .O(doutb[53]),
  .I0(dpb_inst_6_doutb[53]),
  .I1(dpb_inst_7_doutb[53]),
  .S0(dff_q_1)
);
MUX2 mux_inst_182 (
  .O(doutb[54]),
  .I0(dpb_inst_6_doutb[54]),
  .I1(dpb_inst_7_doutb[54]),
  .S0(dff_q_1)
);
MUX2 mux_inst_183 (
  .O(doutb[55]),
  .I0(dpb_inst_6_doutb[55]),
  .I1(dpb_inst_7_doutb[55]),
  .S0(dff_q_1)
);
MUX2 mux_inst_184 (
  .O(doutb[56]),
  .I0(dpb_inst_6_doutb[56]),
  .I1(dpb_inst_7_doutb[56]),
  .S0(dff_q_1)
);
MUX2 mux_inst_185 (
  .O(doutb[57]),
  .I0(dpb_inst_6_doutb[57]),
  .I1(dpb_inst_7_doutb[57]),
  .S0(dff_q_1)
);
MUX2 mux_inst_186 (
  .O(doutb[58]),
  .I0(dpb_inst_6_doutb[58]),
  .I1(dpb_inst_7_doutb[58]),
  .S0(dff_q_1)
);
MUX2 mux_inst_187 (
  .O(doutb[59]),
  .I0(dpb_inst_6_doutb[59]),
  .I1(dpb_inst_7_doutb[59]),
  .S0(dff_q_1)
);
MUX2 mux_inst_188 (
  .O(doutb[60]),
  .I0(dpb_inst_6_doutb[60]),
  .I1(dpb_inst_7_doutb[60]),
  .S0(dff_q_1)
);
MUX2 mux_inst_189 (
  .O(doutb[61]),
  .I0(dpb_inst_6_doutb[61]),
  .I1(dpb_inst_7_doutb[61]),
  .S0(dff_q_1)
);
MUX2 mux_inst_190 (
  .O(doutb[62]),
  .I0(dpb_inst_6_doutb[62]),
  .I1(dpb_inst_7_doutb[62]),
  .S0(dff_q_1)
);
MUX2 mux_inst_191 (
  .O(doutb[63]),
  .I0(dpb_inst_6_doutb[63]),
  .I1(dpb_inst_7_doutb[63]),
  .S0(dff_q_1)
);
MUX2 mux_inst_192 (
  .O(doutb[64]),
  .I0(dpb_inst_8_doutb[64]),
  .I1(dpb_inst_9_doutb[64]),
  .S0(dff_q_1)
);
MUX2 mux_inst_193 (
  .O(doutb[65]),
  .I0(dpb_inst_8_doutb[65]),
  .I1(dpb_inst_9_doutb[65]),
  .S0(dff_q_1)
);
MUX2 mux_inst_194 (
  .O(doutb[66]),
  .I0(dpb_inst_8_doutb[66]),
  .I1(dpb_inst_9_doutb[66]),
  .S0(dff_q_1)
);
MUX2 mux_inst_195 (
  .O(doutb[67]),
  .I0(dpb_inst_8_doutb[67]),
  .I1(dpb_inst_9_doutb[67]),
  .S0(dff_q_1)
);
MUX2 mux_inst_196 (
  .O(doutb[68]),
  .I0(dpb_inst_8_doutb[68]),
  .I1(dpb_inst_9_doutb[68]),
  .S0(dff_q_1)
);
MUX2 mux_inst_197 (
  .O(doutb[69]),
  .I0(dpb_inst_8_doutb[69]),
  .I1(dpb_inst_9_doutb[69]),
  .S0(dff_q_1)
);
MUX2 mux_inst_198 (
  .O(doutb[70]),
  .I0(dpb_inst_8_doutb[70]),
  .I1(dpb_inst_9_doutb[70]),
  .S0(dff_q_1)
);
MUX2 mux_inst_199 (
  .O(doutb[71]),
  .I0(dpb_inst_8_doutb[71]),
  .I1(dpb_inst_9_doutb[71]),
  .S0(dff_q_1)
);
MUX2 mux_inst_200 (
  .O(doutb[72]),
  .I0(dpb_inst_8_doutb[72]),
  .I1(dpb_inst_9_doutb[72]),
  .S0(dff_q_1)
);
MUX2 mux_inst_201 (
  .O(doutb[73]),
  .I0(dpb_inst_8_doutb[73]),
  .I1(dpb_inst_9_doutb[73]),
  .S0(dff_q_1)
);
MUX2 mux_inst_202 (
  .O(doutb[74]),
  .I0(dpb_inst_8_doutb[74]),
  .I1(dpb_inst_9_doutb[74]),
  .S0(dff_q_1)
);
MUX2 mux_inst_203 (
  .O(doutb[75]),
  .I0(dpb_inst_8_doutb[75]),
  .I1(dpb_inst_9_doutb[75]),
  .S0(dff_q_1)
);
MUX2 mux_inst_204 (
  .O(doutb[76]),
  .I0(dpb_inst_8_doutb[76]),
  .I1(dpb_inst_9_doutb[76]),
  .S0(dff_q_1)
);
MUX2 mux_inst_205 (
  .O(doutb[77]),
  .I0(dpb_inst_8_doutb[77]),
  .I1(dpb_inst_9_doutb[77]),
  .S0(dff_q_1)
);
MUX2 mux_inst_206 (
  .O(doutb[78]),
  .I0(dpb_inst_8_doutb[78]),
  .I1(dpb_inst_9_doutb[78]),
  .S0(dff_q_1)
);
MUX2 mux_inst_207 (
  .O(doutb[79]),
  .I0(dpb_inst_8_doutb[79]),
  .I1(dpb_inst_9_doutb[79]),
  .S0(dff_q_1)
);
MUX2 mux_inst_208 (
  .O(doutb[80]),
  .I0(dpb_inst_10_doutb[80]),
  .I1(dpb_inst_11_doutb[80]),
  .S0(dff_q_1)
);
MUX2 mux_inst_209 (
  .O(doutb[81]),
  .I0(dpb_inst_10_doutb[81]),
  .I1(dpb_inst_11_doutb[81]),
  .S0(dff_q_1)
);
MUX2 mux_inst_210 (
  .O(doutb[82]),
  .I0(dpb_inst_10_doutb[82]),
  .I1(dpb_inst_11_doutb[82]),
  .S0(dff_q_1)
);
MUX2 mux_inst_211 (
  .O(doutb[83]),
  .I0(dpb_inst_10_doutb[83]),
  .I1(dpb_inst_11_doutb[83]),
  .S0(dff_q_1)
);
MUX2 mux_inst_212 (
  .O(doutb[84]),
  .I0(dpb_inst_10_doutb[84]),
  .I1(dpb_inst_11_doutb[84]),
  .S0(dff_q_1)
);
MUX2 mux_inst_213 (
  .O(doutb[85]),
  .I0(dpb_inst_10_doutb[85]),
  .I1(dpb_inst_11_doutb[85]),
  .S0(dff_q_1)
);
MUX2 mux_inst_214 (
  .O(doutb[86]),
  .I0(dpb_inst_10_doutb[86]),
  .I1(dpb_inst_11_doutb[86]),
  .S0(dff_q_1)
);
MUX2 mux_inst_215 (
  .O(doutb[87]),
  .I0(dpb_inst_10_doutb[87]),
  .I1(dpb_inst_11_doutb[87]),
  .S0(dff_q_1)
);
MUX2 mux_inst_216 (
  .O(doutb[88]),
  .I0(dpb_inst_10_doutb[88]),
  .I1(dpb_inst_11_doutb[88]),
  .S0(dff_q_1)
);
MUX2 mux_inst_217 (
  .O(doutb[89]),
  .I0(dpb_inst_10_doutb[89]),
  .I1(dpb_inst_11_doutb[89]),
  .S0(dff_q_1)
);
MUX2 mux_inst_218 (
  .O(doutb[90]),
  .I0(dpb_inst_10_doutb[90]),
  .I1(dpb_inst_11_doutb[90]),
  .S0(dff_q_1)
);
MUX2 mux_inst_219 (
  .O(doutb[91]),
  .I0(dpb_inst_10_doutb[91]),
  .I1(dpb_inst_11_doutb[91]),
  .S0(dff_q_1)
);
MUX2 mux_inst_220 (
  .O(doutb[92]),
  .I0(dpb_inst_10_doutb[92]),
  .I1(dpb_inst_11_doutb[92]),
  .S0(dff_q_1)
);
MUX2 mux_inst_221 (
  .O(doutb[93]),
  .I0(dpb_inst_10_doutb[93]),
  .I1(dpb_inst_11_doutb[93]),
  .S0(dff_q_1)
);
MUX2 mux_inst_222 (
  .O(doutb[94]),
  .I0(dpb_inst_10_doutb[94]),
  .I1(dpb_inst_11_doutb[94]),
  .S0(dff_q_1)
);
MUX2 mux_inst_223 (
  .O(doutb[95]),
  .I0(dpb_inst_10_doutb[95]),
  .I1(dpb_inst_11_doutb[95]),
  .S0(dff_q_1)
);
MUX2 mux_inst_224 (
  .O(doutb[96]),
  .I0(dpb_inst_12_doutb[96]),
  .I1(dpb_inst_13_doutb[96]),
  .S0(dff_q_1)
);
MUX2 mux_inst_225 (
  .O(doutb[97]),
  .I0(dpb_inst_12_doutb[97]),
  .I1(dpb_inst_13_doutb[97]),
  .S0(dff_q_1)
);
MUX2 mux_inst_226 (
  .O(doutb[98]),
  .I0(dpb_inst_12_doutb[98]),
  .I1(dpb_inst_13_doutb[98]),
  .S0(dff_q_1)
);
MUX2 mux_inst_227 (
  .O(doutb[99]),
  .I0(dpb_inst_12_doutb[99]),
  .I1(dpb_inst_13_doutb[99]),
  .S0(dff_q_1)
);
MUX2 mux_inst_228 (
  .O(doutb[100]),
  .I0(dpb_inst_12_doutb[100]),
  .I1(dpb_inst_13_doutb[100]),
  .S0(dff_q_1)
);
MUX2 mux_inst_229 (
  .O(doutb[101]),
  .I0(dpb_inst_12_doutb[101]),
  .I1(dpb_inst_13_doutb[101]),
  .S0(dff_q_1)
);
MUX2 mux_inst_230 (
  .O(doutb[102]),
  .I0(dpb_inst_12_doutb[102]),
  .I1(dpb_inst_13_doutb[102]),
  .S0(dff_q_1)
);
MUX2 mux_inst_231 (
  .O(doutb[103]),
  .I0(dpb_inst_12_doutb[103]),
  .I1(dpb_inst_13_doutb[103]),
  .S0(dff_q_1)
);
MUX2 mux_inst_232 (
  .O(doutb[104]),
  .I0(dpb_inst_12_doutb[104]),
  .I1(dpb_inst_13_doutb[104]),
  .S0(dff_q_1)
);
MUX2 mux_inst_233 (
  .O(doutb[105]),
  .I0(dpb_inst_12_doutb[105]),
  .I1(dpb_inst_13_doutb[105]),
  .S0(dff_q_1)
);
MUX2 mux_inst_234 (
  .O(doutb[106]),
  .I0(dpb_inst_12_doutb[106]),
  .I1(dpb_inst_13_doutb[106]),
  .S0(dff_q_1)
);
MUX2 mux_inst_235 (
  .O(doutb[107]),
  .I0(dpb_inst_12_doutb[107]),
  .I1(dpb_inst_13_doutb[107]),
  .S0(dff_q_1)
);
MUX2 mux_inst_236 (
  .O(doutb[108]),
  .I0(dpb_inst_12_doutb[108]),
  .I1(dpb_inst_13_doutb[108]),
  .S0(dff_q_1)
);
MUX2 mux_inst_237 (
  .O(doutb[109]),
  .I0(dpb_inst_12_doutb[109]),
  .I1(dpb_inst_13_doutb[109]),
  .S0(dff_q_1)
);
MUX2 mux_inst_238 (
  .O(doutb[110]),
  .I0(dpb_inst_12_doutb[110]),
  .I1(dpb_inst_13_doutb[110]),
  .S0(dff_q_1)
);
MUX2 mux_inst_239 (
  .O(doutb[111]),
  .I0(dpb_inst_12_doutb[111]),
  .I1(dpb_inst_13_doutb[111]),
  .S0(dff_q_1)
);
MUX2 mux_inst_240 (
  .O(doutb[112]),
  .I0(dpb_inst_14_doutb[112]),
  .I1(dpb_inst_15_doutb[112]),
  .S0(dff_q_1)
);
MUX2 mux_inst_241 (
  .O(doutb[113]),
  .I0(dpb_inst_14_doutb[113]),
  .I1(dpb_inst_15_doutb[113]),
  .S0(dff_q_1)
);
MUX2 mux_inst_242 (
  .O(doutb[114]),
  .I0(dpb_inst_14_doutb[114]),
  .I1(dpb_inst_15_doutb[114]),
  .S0(dff_q_1)
);
MUX2 mux_inst_243 (
  .O(doutb[115]),
  .I0(dpb_inst_14_doutb[115]),
  .I1(dpb_inst_15_doutb[115]),
  .S0(dff_q_1)
);
MUX2 mux_inst_244 (
  .O(doutb[116]),
  .I0(dpb_inst_14_doutb[116]),
  .I1(dpb_inst_15_doutb[116]),
  .S0(dff_q_1)
);
MUX2 mux_inst_245 (
  .O(doutb[117]),
  .I0(dpb_inst_14_doutb[117]),
  .I1(dpb_inst_15_doutb[117]),
  .S0(dff_q_1)
);
MUX2 mux_inst_246 (
  .O(doutb[118]),
  .I0(dpb_inst_14_doutb[118]),
  .I1(dpb_inst_15_doutb[118]),
  .S0(dff_q_1)
);
MUX2 mux_inst_247 (
  .O(doutb[119]),
  .I0(dpb_inst_14_doutb[119]),
  .I1(dpb_inst_15_doutb[119]),
  .S0(dff_q_1)
);
MUX2 mux_inst_248 (
  .O(doutb[120]),
  .I0(dpb_inst_14_doutb[120]),
  .I1(dpb_inst_15_doutb[120]),
  .S0(dff_q_1)
);
MUX2 mux_inst_249 (
  .O(doutb[121]),
  .I0(dpb_inst_14_doutb[121]),
  .I1(dpb_inst_15_doutb[121]),
  .S0(dff_q_1)
);
MUX2 mux_inst_250 (
  .O(doutb[122]),
  .I0(dpb_inst_14_doutb[122]),
  .I1(dpb_inst_15_doutb[122]),
  .S0(dff_q_1)
);
MUX2 mux_inst_251 (
  .O(doutb[123]),
  .I0(dpb_inst_14_doutb[123]),
  .I1(dpb_inst_15_doutb[123]),
  .S0(dff_q_1)
);
MUX2 mux_inst_252 (
  .O(doutb[124]),
  .I0(dpb_inst_14_doutb[124]),
  .I1(dpb_inst_15_doutb[124]),
  .S0(dff_q_1)
);
MUX2 mux_inst_253 (
  .O(doutb[125]),
  .I0(dpb_inst_14_doutb[125]),
  .I1(dpb_inst_15_doutb[125]),
  .S0(dff_q_1)
);
MUX2 mux_inst_254 (
  .O(doutb[126]),
  .I0(dpb_inst_14_doutb[126]),
  .I1(dpb_inst_15_doutb[126]),
  .S0(dff_q_1)
);
MUX2 mux_inst_255 (
  .O(doutb[127]),
  .I0(dpb_inst_14_doutb[127]),
  .I1(dpb_inst_15_doutb[127]),
  .S0(dff_q_1)
);
endmodule //Gowin_DPB_128_2048
