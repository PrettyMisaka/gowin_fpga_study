module ddr3_master_cmd(

);

endmodule