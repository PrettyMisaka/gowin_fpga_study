module sdio_init(
    input clk48mhz,
    input rst_n,

    input   sdio_cmd_i  ,
    output  reg sdio_cmd_o  ,
    output  reg sdio_cmd_oen,

    output wire sdio_clk,

    output  reg init_down
);



endmodule